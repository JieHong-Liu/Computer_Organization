module Control
(
    input Run,
    input Reset,
    input clk,
    input LSB,
    output W_ctrl,
    output [5:0]ADDU_ctrl,
    output SRL_ctrl,
    output Ready
);


endmodule
