module Multiplicand(Reset,W_ctrl,Multiplicand_in,Multiplicand_out);
    input Reset;
    input W_ctrl;
    input [31:0]Multiplicand_in;
    output [31:0]Multiplicand_out;
endmodule
