module CompMultiplier(
    input clk,
    input Reset,
    input Run,
    input [31:0] Multiplier_in,
    input [31:0] Multiplicand_in,
    output [63:0]Product_out,
    output Ready
);
endmodule
