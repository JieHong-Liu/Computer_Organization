module ALU(
    input   [31:0]  Src1,
    input   [31:0]  Src2,
    input   [4:0]   Shamt,
    input   [5:0]   Funct,
    output  [31:0]  result
);


endmodule