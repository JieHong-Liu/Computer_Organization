module tb_ID_EX(

);



endmodule