module ALU(
    input [31:0]Src1,
    input [31:0]Src2,
    output [31:0]Result,
    output Carry
);
endmodule
