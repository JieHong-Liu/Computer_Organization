module Control(
    input [5:0] OpCode,
    output wire RegWrite
);

endmodule