module Product(
    input SRL_ctrl,
    input W_ctrl,
    input Ready,
    input Reset,
    input clk,
    input ALU_carry,
    input [31:0]ALU_Result,
    input [31:0]Multiplier_in,
    output [63:0]Product_out
);

endmodule
